// nios2_control.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module nios2_control (
		input  wire [3:0] button_pio_external_in_port,            //             button_pio_external.in_port
		output wire [3:0] button_pio_external_out_port,           //                                .out_port
		input  wire       clk_clk,                                //                             clk.clk
		output wire [7:0] led_led_pio_external_connection_export, // led_led_pio_external_connection.export
		input  wire       reset_reset_n                           //                           reset.reset_n
	);

	wire         altpll_0_c0_clk;                                             // altpll_0:c0 -> [altpll_0:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, mm_interconnect_0:altpll_0_c0_clk, nios2_cpu:clk, onchip_flash_0:clock, onchip_ram:clk, rst_controller:clk, slow_periph_bridge:s0_clk]
	wire         altpll_0_c1_clk;                                             // altpll_0:c1 -> [button_pio:clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, irq_synchronizer_002:receiver_clk, jtag_uart_0:clk, led_pio:clk, mm_interconnect_1:altpll_0_c1_clk, rst_controller_001:clk, slow_periph_bridge:m0_clk, sysid:clock, timer_0:clk]
	wire  [31:0] nios2_cpu_data_master_readdata;                              // mm_interconnect_0:nios2_cpu_data_master_readdata -> nios2_cpu:d_readdata
	wire         nios2_cpu_data_master_waitrequest;                           // mm_interconnect_0:nios2_cpu_data_master_waitrequest -> nios2_cpu:d_waitrequest
	wire         nios2_cpu_data_master_debugaccess;                           // nios2_cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_cpu_data_master_debugaccess
	wire  [21:0] nios2_cpu_data_master_address;                               // nios2_cpu:d_address -> mm_interconnect_0:nios2_cpu_data_master_address
	wire   [3:0] nios2_cpu_data_master_byteenable;                            // nios2_cpu:d_byteenable -> mm_interconnect_0:nios2_cpu_data_master_byteenable
	wire         nios2_cpu_data_master_read;                                  // nios2_cpu:d_read -> mm_interconnect_0:nios2_cpu_data_master_read
	wire         nios2_cpu_data_master_readdatavalid;                         // mm_interconnect_0:nios2_cpu_data_master_readdatavalid -> nios2_cpu:d_readdatavalid
	wire         nios2_cpu_data_master_write;                                 // nios2_cpu:d_write -> mm_interconnect_0:nios2_cpu_data_master_write
	wire  [31:0] nios2_cpu_data_master_writedata;                             // nios2_cpu:d_writedata -> mm_interconnect_0:nios2_cpu_data_master_writedata
	wire  [31:0] nios2_cpu_instruction_master_readdata;                       // mm_interconnect_0:nios2_cpu_instruction_master_readdata -> nios2_cpu:i_readdata
	wire         nios2_cpu_instruction_master_waitrequest;                    // mm_interconnect_0:nios2_cpu_instruction_master_waitrequest -> nios2_cpu:i_waitrequest
	wire  [21:0] nios2_cpu_instruction_master_address;                        // nios2_cpu:i_address -> mm_interconnect_0:nios2_cpu_instruction_master_address
	wire         nios2_cpu_instruction_master_read;                           // nios2_cpu:i_read -> mm_interconnect_0:nios2_cpu_instruction_master_read
	wire         nios2_cpu_instruction_master_readdatavalid;                  // mm_interconnect_0:nios2_cpu_instruction_master_readdatavalid -> nios2_cpu:i_readdatavalid
	wire  [31:0] mm_interconnect_0_onchip_flash_0_csr_readdata;               // onchip_flash_0:avmm_csr_readdata -> mm_interconnect_0:onchip_flash_0_csr_readdata
	wire   [0:0] mm_interconnect_0_onchip_flash_0_csr_address;                // mm_interconnect_0:onchip_flash_0_csr_address -> onchip_flash_0:avmm_csr_addr
	wire         mm_interconnect_0_onchip_flash_0_csr_read;                   // mm_interconnect_0:onchip_flash_0_csr_read -> onchip_flash_0:avmm_csr_read
	wire         mm_interconnect_0_onchip_flash_0_csr_write;                  // mm_interconnect_0:onchip_flash_0_csr_write -> onchip_flash_0:avmm_csr_write
	wire  [31:0] mm_interconnect_0_onchip_flash_0_csr_writedata;              // mm_interconnect_0:onchip_flash_0_csr_writedata -> onchip_flash_0:avmm_csr_writedata
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_readdata;              // onchip_flash_0:avmm_data_readdata -> mm_interconnect_0:onchip_flash_0_data_readdata
	wire         mm_interconnect_0_onchip_flash_0_data_waitrequest;           // onchip_flash_0:avmm_data_waitrequest -> mm_interconnect_0:onchip_flash_0_data_waitrequest
	wire  [16:0] mm_interconnect_0_onchip_flash_0_data_address;               // mm_interconnect_0:onchip_flash_0_data_address -> onchip_flash_0:avmm_data_addr
	wire         mm_interconnect_0_onchip_flash_0_data_read;                  // mm_interconnect_0:onchip_flash_0_data_read -> onchip_flash_0:avmm_data_read
	wire         mm_interconnect_0_onchip_flash_0_data_readdatavalid;         // onchip_flash_0:avmm_data_readdatavalid -> mm_interconnect_0:onchip_flash_0_data_readdatavalid
	wire         mm_interconnect_0_onchip_flash_0_data_write;                 // mm_interconnect_0:onchip_flash_0_data_write -> onchip_flash_0:avmm_data_write
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_writedata;             // mm_interconnect_0:onchip_flash_0_data_writedata -> onchip_flash_0:avmm_data_writedata
	wire   [3:0] mm_interconnect_0_onchip_flash_0_data_burstcount;            // mm_interconnect_0:onchip_flash_0_data_burstcount -> onchip_flash_0:avmm_data_burstcount
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata;        // nios2_cpu:debug_mem_slave_readdata -> mm_interconnect_0:nios2_cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest;     // nios2_cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess;     // mm_interconnect_0:nios2_cpu_debug_mem_slave_debugaccess -> nios2_cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_address;         // mm_interconnect_0:nios2_cpu_debug_mem_slave_address -> nios2_cpu:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_read;            // mm_interconnect_0:nios2_cpu_debug_mem_slave_read -> nios2_cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable;      // mm_interconnect_0:nios2_cpu_debug_mem_slave_byteenable -> nios2_cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_write;           // mm_interconnect_0:nios2_cpu_debug_mem_slave_write -> nios2_cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata;       // mm_interconnect_0:nios2_cpu_debug_mem_slave_writedata -> nios2_cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;               // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;                // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                   // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                  // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;              // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire  [31:0] mm_interconnect_0_slow_periph_bridge_s0_readdata;            // slow_periph_bridge:s0_readdata -> mm_interconnect_0:slow_periph_bridge_s0_readdata
	wire         mm_interconnect_0_slow_periph_bridge_s0_waitrequest;         // slow_periph_bridge:s0_waitrequest -> mm_interconnect_0:slow_periph_bridge_s0_waitrequest
	wire         mm_interconnect_0_slow_periph_bridge_s0_debugaccess;         // mm_interconnect_0:slow_periph_bridge_s0_debugaccess -> slow_periph_bridge:s0_debugaccess
	wire   [9:0] mm_interconnect_0_slow_periph_bridge_s0_address;             // mm_interconnect_0:slow_periph_bridge_s0_address -> slow_periph_bridge:s0_address
	wire         mm_interconnect_0_slow_periph_bridge_s0_read;                // mm_interconnect_0:slow_periph_bridge_s0_read -> slow_periph_bridge:s0_read
	wire   [3:0] mm_interconnect_0_slow_periph_bridge_s0_byteenable;          // mm_interconnect_0:slow_periph_bridge_s0_byteenable -> slow_periph_bridge:s0_byteenable
	wire         mm_interconnect_0_slow_periph_bridge_s0_readdatavalid;       // slow_periph_bridge:s0_readdatavalid -> mm_interconnect_0:slow_periph_bridge_s0_readdatavalid
	wire         mm_interconnect_0_slow_periph_bridge_s0_write;               // mm_interconnect_0:slow_periph_bridge_s0_write -> slow_periph_bridge:s0_write
	wire  [31:0] mm_interconnect_0_slow_periph_bridge_s0_writedata;           // mm_interconnect_0:slow_periph_bridge_s0_writedata -> slow_periph_bridge:s0_writedata
	wire   [0:0] mm_interconnect_0_slow_periph_bridge_s0_burstcount;          // mm_interconnect_0:slow_periph_bridge_s0_burstcount -> slow_periph_bridge:s0_burstcount
	wire         mm_interconnect_0_onchip_ram_s1_chipselect;                  // mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_readdata;                    // onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_ram_s1_address;                     // mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	wire   [3:0] mm_interconnect_0_onchip_ram_s1_byteenable;                  // mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	wire         mm_interconnect_0_onchip_ram_s1_write;                       // mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_writedata;                   // mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	wire         mm_interconnect_0_onchip_ram_s1_clken;                       // mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	wire         slow_periph_bridge_m0_waitrequest;                           // mm_interconnect_1:slow_periph_bridge_m0_waitrequest -> slow_periph_bridge:m0_waitrequest
	wire  [31:0] slow_periph_bridge_m0_readdata;                              // mm_interconnect_1:slow_periph_bridge_m0_readdata -> slow_periph_bridge:m0_readdata
	wire         slow_periph_bridge_m0_debugaccess;                           // slow_periph_bridge:m0_debugaccess -> mm_interconnect_1:slow_periph_bridge_m0_debugaccess
	wire   [9:0] slow_periph_bridge_m0_address;                               // slow_periph_bridge:m0_address -> mm_interconnect_1:slow_periph_bridge_m0_address
	wire         slow_periph_bridge_m0_read;                                  // slow_periph_bridge:m0_read -> mm_interconnect_1:slow_periph_bridge_m0_read
	wire   [3:0] slow_periph_bridge_m0_byteenable;                            // slow_periph_bridge:m0_byteenable -> mm_interconnect_1:slow_periph_bridge_m0_byteenable
	wire         slow_periph_bridge_m0_readdatavalid;                         // mm_interconnect_1:slow_periph_bridge_m0_readdatavalid -> slow_periph_bridge:m0_readdatavalid
	wire  [31:0] slow_periph_bridge_m0_writedata;                             // slow_periph_bridge:m0_writedata -> mm_interconnect_1:slow_periph_bridge_m0_writedata
	wire         slow_periph_bridge_m0_write;                                 // slow_periph_bridge:m0_write -> mm_interconnect_1:slow_periph_bridge_m0_write
	wire   [0:0] slow_periph_bridge_m0_burstcount;                            // slow_periph_bridge:m0_burstcount -> mm_interconnect_1:slow_periph_bridge_m0_burstcount
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;              // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;               // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire         mm_interconnect_1_led_pio_s1_chipselect;                     // mm_interconnect_1:led_pio_s1_chipselect -> led_pio:chipselect
	wire  [31:0] mm_interconnect_1_led_pio_s1_readdata;                       // led_pio:readdata -> mm_interconnect_1:led_pio_s1_readdata
	wire   [1:0] mm_interconnect_1_led_pio_s1_address;                        // mm_interconnect_1:led_pio_s1_address -> led_pio:address
	wire         mm_interconnect_1_led_pio_s1_write;                          // mm_interconnect_1:led_pio_s1_write -> led_pio:write_n
	wire  [31:0] mm_interconnect_1_led_pio_s1_writedata;                      // mm_interconnect_1:led_pio_s1_writedata -> led_pio:writedata
	wire         mm_interconnect_1_button_pio_s1_chipselect;                  // mm_interconnect_1:button_pio_s1_chipselect -> button_pio:chipselect
	wire  [31:0] mm_interconnect_1_button_pio_s1_readdata;                    // button_pio:readdata -> mm_interconnect_1:button_pio_s1_readdata
	wire   [1:0] mm_interconnect_1_button_pio_s1_address;                     // mm_interconnect_1:button_pio_s1_address -> button_pio:address
	wire         mm_interconnect_1_button_pio_s1_write;                       // mm_interconnect_1:button_pio_s1_write -> button_pio:write_n
	wire  [31:0] mm_interconnect_1_button_pio_s1_writedata;                   // mm_interconnect_1:button_pio_s1_writedata -> button_pio:writedata
	wire         mm_interconnect_1_timer_0_s1_chipselect;                     // mm_interconnect_1:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_1_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_1:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_1_timer_0_s1_address;                        // mm_interconnect_1:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_1_timer_0_s1_write;                          // mm_interconnect_1:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_1_timer_0_s1_writedata;                      // mm_interconnect_1:timer_0_s1_writedata -> timer_0:writedata
	wire  [31:0] nios2_cpu_irq_irq;                                           // irq_mapper:sender_irq -> nios2_cpu:irq
	wire         irq_mapper_receiver0_irq;                                    // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                               // button_pio:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                    // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                           // timer_0:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver2_irq;                                    // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                           // jtag_uart_0:av_irq -> irq_synchronizer_002:receiver_irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [altpll_0:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, mm_interconnect_0:nios2_cpu_reset_reset_bridge_in_reset_reset, nios2_cpu:reset_n, onchip_flash_0:reset_n, onchip_ram:reset, rst_translator:in_reset, slow_periph_bridge:s0_reset]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2_cpu:reset_req, onchip_ram:reset_req, rst_translator:reset_req_in]
	wire         nios2_cpu_debug_reset_request_reset;                         // nios2_cpu:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [button_pio:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, jtag_uart_0:rst_n, led_pio:reset_n, mm_interconnect_1:slow_periph_bridge_m0_reset_reset_bridge_in_reset_reset, slow_periph_bridge:m0_reset, sysid:reset_n, timer_0:reset_n]

	nios2_control_altpll_0 altpll_0 (
		.clk                (altpll_0_c0_clk),                                //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                 // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_0_c0_clk),                                //                    c0.clk
		.c1                 (altpll_0_c1_clk),                                //                    c1.clk
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.c2                 (),                                               //           (terminated)
		.c3                 (),                                               //           (terminated)
		.c4                 (),                                               //           (terminated)
		.areset             (1'b0),                                           //           (terminated)
		.locked             (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (3'b000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	nios2_control_button_pio button_pio (
		.clk        (altpll_0_c1_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_1_button_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_button_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_button_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_button_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_button_pio_s1_readdata),   //                    .readdata
		.in_port    (button_pio_external_in_port),                // external_connection.export
		.out_port   (button_pio_external_out_port),               //                    .export
		.irq        (irq_synchronizer_receiver_irq)               //                 irq.irq
	);

	nios2_control_jtag_uart_0 jtag_uart_0 (
		.clk            (altpll_0_c1_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_002_receiver_irq)                            //               irq.irq
	);

	nios2_control_led_pio led_pio (
		.clk        (altpll_0_c1_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_pio_s1_readdata),   //                    .readdata
		.out_port   (led_led_pio_external_connection_export)   // external_connection.export
	);

	nios2_control_nios2_cpu nios2_cpu (
		.clk                                 (altpll_0_c0_clk),                                         //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                         //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                      //                          .reset_req
		.d_address                           (nios2_cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_cpu_data_master_read),                              //                          .read
		.d_readdata                          (nios2_cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_cpu_data_master_write),                             //                          .write
		.d_writedata                         (nios2_cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                         // custom_instruction_master.readra
	);

	altera_onchip_flash #(
		.INIT_FILENAME                       (""),
		.INIT_FILENAME_SIM                   (""),
		.DEVICE_FAMILY                       ("MAX 10"),
		.PART_NAME                           ("10M08DAF484C8GES"),
		.DEVICE_ID                           ("08"),
		.SECTOR1_START_ADDR                  (0),
		.SECTOR1_END_ADDR                    (4095),
		.SECTOR2_START_ADDR                  (4096),
		.SECTOR2_END_ADDR                    (8191),
		.SECTOR3_START_ADDR                  (8192),
		.SECTOR3_END_ADDR                    (29183),
		.SECTOR4_START_ADDR                  (29184),
		.SECTOR4_END_ADDR                    (44031),
		.SECTOR5_START_ADDR                  (44032),
		.SECTOR5_END_ADDR                    (79871),
		.MIN_VALID_ADDR                      (0),
		.MAX_VALID_ADDR                      (79871),
		.MIN_UFM_VALID_ADDR                  (0),
		.MAX_UFM_VALID_ADDR                  (29183),
		.SECTOR1_MAP                         (1),
		.SECTOR2_MAP                         (2),
		.SECTOR3_MAP                         (3),
		.SECTOR4_MAP                         (4),
		.SECTOR5_MAP                         (5),
		.ADDR_RANGE1_END_ADDR                (79871),
		.ADDR_RANGE1_OFFSET                  (512),
		.ADDR_RANGE2_OFFSET                  (0),
		.AVMM_DATA_ADDR_WIDTH                (17),
		.AVMM_DATA_DATA_WIDTH                (32),
		.AVMM_DATA_BURSTCOUNT_WIDTH          (4),
		.SECTOR_READ_PROTECTION_MODE         (4),
		.FLASH_SEQ_READ_DATA_COUNT           (2),
		.FLASH_ADDR_ALIGNMENT_BITS           (1),
		.FLASH_READ_CYCLE_MAX_INDEX          (4),
		.FLASH_RESET_CYCLE_MAX_INDEX         (20),
		.FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  (96),
		.FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX (28000000),
		.FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX (24400),
		.PARALLEL_MODE                       (1),
		.READ_AND_WRITE_MODE                 (1),
		.WRAPPING_BURST_MODE                 (0),
		.IS_DUAL_BOOT                        ("False"),
		.IS_ERAM_SKIP                        ("True"),
		.IS_COMPRESSED_IMAGE                 ("False")
	) onchip_flash_0 (
		.clock                   (altpll_0_c0_clk),                                     //    clk.clk
		.reset_n                 (~rst_controller_reset_out_reset),                     // nreset.reset_n
		.avmm_data_addr          (mm_interconnect_0_onchip_flash_0_data_address),       //   data.address
		.avmm_data_read          (mm_interconnect_0_onchip_flash_0_data_read),          //       .read
		.avmm_data_writedata     (mm_interconnect_0_onchip_flash_0_data_writedata),     //       .writedata
		.avmm_data_write         (mm_interconnect_0_onchip_flash_0_data_write),         //       .write
		.avmm_data_readdata      (mm_interconnect_0_onchip_flash_0_data_readdata),      //       .readdata
		.avmm_data_waitrequest   (mm_interconnect_0_onchip_flash_0_data_waitrequest),   //       .waitrequest
		.avmm_data_readdatavalid (mm_interconnect_0_onchip_flash_0_data_readdatavalid), //       .readdatavalid
		.avmm_data_burstcount    (mm_interconnect_0_onchip_flash_0_data_burstcount),    //       .burstcount
		.avmm_csr_addr           (mm_interconnect_0_onchip_flash_0_csr_address),        //    csr.address
		.avmm_csr_read           (mm_interconnect_0_onchip_flash_0_csr_read),           //       .read
		.avmm_csr_writedata      (mm_interconnect_0_onchip_flash_0_csr_writedata),      //       .writedata
		.avmm_csr_write          (mm_interconnect_0_onchip_flash_0_csr_write),          //       .write
		.avmm_csr_readdata       (mm_interconnect_0_onchip_flash_0_csr_readdata)        //       .readdata
	);

	nios2_control_onchip_ram onchip_ram (
		.clk        (altpll_0_c0_clk),                            //   clk1.clk
		.address    (mm_interconnect_0_onchip_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                        // (terminated)
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (32),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) slow_periph_bridge (
		.m0_clk           (altpll_0_c1_clk),                                       //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                    // m0_reset.reset
		.s0_clk           (altpll_0_c0_clk),                                       //   s0_clk.clk
		.s0_reset         (rst_controller_reset_out_reset),                        // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_slow_periph_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_slow_periph_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_slow_periph_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_slow_periph_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_slow_periph_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_slow_periph_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_slow_periph_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_slow_periph_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_slow_periph_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_slow_periph_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (slow_periph_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (slow_periph_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (slow_periph_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (slow_periph_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (slow_periph_bridge_m0_writedata),                       //         .writedata
		.m0_address       (slow_periph_bridge_m0_address),                         //         .address
		.m0_write         (slow_periph_bridge_m0_write),                           //         .write
		.m0_read          (slow_periph_bridge_m0_read),                            //         .read
		.m0_byteenable    (slow_periph_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (slow_periph_bridge_m0_debugaccess)                      //         .debugaccess
	);

	nios2_control_sysid sysid (
		.clock    (altpll_0_c1_clk),                                //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	nios2_control_timer_0 timer_0 (
		.clk        (altpll_0_c1_clk),                         //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_1_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_0_s1_write),     //      .write_n
		.irq        (irq_synchronizer_001_receiver_irq)        //   irq.irq
	);

	nios2_control_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                             (altpll_0_c0_clk),                                         //                           altpll_0_c0.clk
		.nios2_cpu_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                          // nios2_cpu_reset_reset_bridge_in_reset.reset
		.nios2_cpu_data_master_address               (nios2_cpu_data_master_address),                           //                 nios2_cpu_data_master.address
		.nios2_cpu_data_master_waitrequest           (nios2_cpu_data_master_waitrequest),                       //                                      .waitrequest
		.nios2_cpu_data_master_byteenable            (nios2_cpu_data_master_byteenable),                        //                                      .byteenable
		.nios2_cpu_data_master_read                  (nios2_cpu_data_master_read),                              //                                      .read
		.nios2_cpu_data_master_readdata              (nios2_cpu_data_master_readdata),                          //                                      .readdata
		.nios2_cpu_data_master_readdatavalid         (nios2_cpu_data_master_readdatavalid),                     //                                      .readdatavalid
		.nios2_cpu_data_master_write                 (nios2_cpu_data_master_write),                             //                                      .write
		.nios2_cpu_data_master_writedata             (nios2_cpu_data_master_writedata),                         //                                      .writedata
		.nios2_cpu_data_master_debugaccess           (nios2_cpu_data_master_debugaccess),                       //                                      .debugaccess
		.nios2_cpu_instruction_master_address        (nios2_cpu_instruction_master_address),                    //          nios2_cpu_instruction_master.address
		.nios2_cpu_instruction_master_waitrequest    (nios2_cpu_instruction_master_waitrequest),                //                                      .waitrequest
		.nios2_cpu_instruction_master_read           (nios2_cpu_instruction_master_read),                       //                                      .read
		.nios2_cpu_instruction_master_readdata       (nios2_cpu_instruction_master_readdata),                   //                                      .readdata
		.nios2_cpu_instruction_master_readdatavalid  (nios2_cpu_instruction_master_readdatavalid),              //                                      .readdatavalid
		.altpll_0_pll_slave_address                  (mm_interconnect_0_altpll_0_pll_slave_address),            //                    altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                    (mm_interconnect_0_altpll_0_pll_slave_write),              //                                      .write
		.altpll_0_pll_slave_read                     (mm_interconnect_0_altpll_0_pll_slave_read),               //                                      .read
		.altpll_0_pll_slave_readdata                 (mm_interconnect_0_altpll_0_pll_slave_readdata),           //                                      .readdata
		.altpll_0_pll_slave_writedata                (mm_interconnect_0_altpll_0_pll_slave_writedata),          //                                      .writedata
		.nios2_cpu_debug_mem_slave_address           (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),     //             nios2_cpu_debug_mem_slave.address
		.nios2_cpu_debug_mem_slave_write             (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),       //                                      .write
		.nios2_cpu_debug_mem_slave_read              (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),        //                                      .read
		.nios2_cpu_debug_mem_slave_readdata          (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),    //                                      .readdata
		.nios2_cpu_debug_mem_slave_writedata         (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),   //                                      .writedata
		.nios2_cpu_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),  //                                      .byteenable
		.nios2_cpu_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest), //                                      .waitrequest
		.nios2_cpu_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess), //                                      .debugaccess
		.onchip_flash_0_csr_address                  (mm_interconnect_0_onchip_flash_0_csr_address),            //                    onchip_flash_0_csr.address
		.onchip_flash_0_csr_write                    (mm_interconnect_0_onchip_flash_0_csr_write),              //                                      .write
		.onchip_flash_0_csr_read                     (mm_interconnect_0_onchip_flash_0_csr_read),               //                                      .read
		.onchip_flash_0_csr_readdata                 (mm_interconnect_0_onchip_flash_0_csr_readdata),           //                                      .readdata
		.onchip_flash_0_csr_writedata                (mm_interconnect_0_onchip_flash_0_csr_writedata),          //                                      .writedata
		.onchip_flash_0_data_address                 (mm_interconnect_0_onchip_flash_0_data_address),           //                   onchip_flash_0_data.address
		.onchip_flash_0_data_write                   (mm_interconnect_0_onchip_flash_0_data_write),             //                                      .write
		.onchip_flash_0_data_read                    (mm_interconnect_0_onchip_flash_0_data_read),              //                                      .read
		.onchip_flash_0_data_readdata                (mm_interconnect_0_onchip_flash_0_data_readdata),          //                                      .readdata
		.onchip_flash_0_data_writedata               (mm_interconnect_0_onchip_flash_0_data_writedata),         //                                      .writedata
		.onchip_flash_0_data_burstcount              (mm_interconnect_0_onchip_flash_0_data_burstcount),        //                                      .burstcount
		.onchip_flash_0_data_readdatavalid           (mm_interconnect_0_onchip_flash_0_data_readdatavalid),     //                                      .readdatavalid
		.onchip_flash_0_data_waitrequest             (mm_interconnect_0_onchip_flash_0_data_waitrequest),       //                                      .waitrequest
		.onchip_ram_s1_address                       (mm_interconnect_0_onchip_ram_s1_address),                 //                         onchip_ram_s1.address
		.onchip_ram_s1_write                         (mm_interconnect_0_onchip_ram_s1_write),                   //                                      .write
		.onchip_ram_s1_readdata                      (mm_interconnect_0_onchip_ram_s1_readdata),                //                                      .readdata
		.onchip_ram_s1_writedata                     (mm_interconnect_0_onchip_ram_s1_writedata),               //                                      .writedata
		.onchip_ram_s1_byteenable                    (mm_interconnect_0_onchip_ram_s1_byteenable),              //                                      .byteenable
		.onchip_ram_s1_chipselect                    (mm_interconnect_0_onchip_ram_s1_chipselect),              //                                      .chipselect
		.onchip_ram_s1_clken                         (mm_interconnect_0_onchip_ram_s1_clken),                   //                                      .clken
		.slow_periph_bridge_s0_address               (mm_interconnect_0_slow_periph_bridge_s0_address),         //                 slow_periph_bridge_s0.address
		.slow_periph_bridge_s0_write                 (mm_interconnect_0_slow_periph_bridge_s0_write),           //                                      .write
		.slow_periph_bridge_s0_read                  (mm_interconnect_0_slow_periph_bridge_s0_read),            //                                      .read
		.slow_periph_bridge_s0_readdata              (mm_interconnect_0_slow_periph_bridge_s0_readdata),        //                                      .readdata
		.slow_periph_bridge_s0_writedata             (mm_interconnect_0_slow_periph_bridge_s0_writedata),       //                                      .writedata
		.slow_periph_bridge_s0_burstcount            (mm_interconnect_0_slow_periph_bridge_s0_burstcount),      //                                      .burstcount
		.slow_periph_bridge_s0_byteenable            (mm_interconnect_0_slow_periph_bridge_s0_byteenable),      //                                      .byteenable
		.slow_periph_bridge_s0_readdatavalid         (mm_interconnect_0_slow_periph_bridge_s0_readdatavalid),   //                                      .readdatavalid
		.slow_periph_bridge_s0_waitrequest           (mm_interconnect_0_slow_periph_bridge_s0_waitrequest),     //                                      .waitrequest
		.slow_periph_bridge_s0_debugaccess           (mm_interconnect_0_slow_periph_bridge_s0_debugaccess)      //                                      .debugaccess
	);

	nios2_control_mm_interconnect_1 mm_interconnect_1 (
		.altpll_0_c1_clk                                         (altpll_0_c1_clk),                                             //                                       altpll_0_c1.clk
		.slow_periph_bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // slow_periph_bridge_m0_reset_reset_bridge_in_reset.reset
		.slow_periph_bridge_m0_address                           (slow_periph_bridge_m0_address),                               //                             slow_periph_bridge_m0.address
		.slow_periph_bridge_m0_waitrequest                       (slow_periph_bridge_m0_waitrequest),                           //                                                  .waitrequest
		.slow_periph_bridge_m0_burstcount                        (slow_periph_bridge_m0_burstcount),                            //                                                  .burstcount
		.slow_periph_bridge_m0_byteenable                        (slow_periph_bridge_m0_byteenable),                            //                                                  .byteenable
		.slow_periph_bridge_m0_read                              (slow_periph_bridge_m0_read),                                  //                                                  .read
		.slow_periph_bridge_m0_readdata                          (slow_periph_bridge_m0_readdata),                              //                                                  .readdata
		.slow_periph_bridge_m0_readdatavalid                     (slow_periph_bridge_m0_readdatavalid),                         //                                                  .readdatavalid
		.slow_periph_bridge_m0_write                             (slow_periph_bridge_m0_write),                                 //                                                  .write
		.slow_periph_bridge_m0_writedata                         (slow_periph_bridge_m0_writedata),                             //                                                  .writedata
		.slow_periph_bridge_m0_debugaccess                       (slow_periph_bridge_m0_debugaccess),                           //                                                  .debugaccess
		.button_pio_s1_address                                   (mm_interconnect_1_button_pio_s1_address),                     //                                     button_pio_s1.address
		.button_pio_s1_write                                     (mm_interconnect_1_button_pio_s1_write),                       //                                                  .write
		.button_pio_s1_readdata                                  (mm_interconnect_1_button_pio_s1_readdata),                    //                                                  .readdata
		.button_pio_s1_writedata                                 (mm_interconnect_1_button_pio_s1_writedata),                   //                                                  .writedata
		.button_pio_s1_chipselect                                (mm_interconnect_1_button_pio_s1_chipselect),                  //                                                  .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                   (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address),     //                     jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                     (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write),       //                                                  .write
		.jtag_uart_0_avalon_jtag_slave_read                      (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read),        //                                                  .read
		.jtag_uart_0_avalon_jtag_slave_readdata                  (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata),    //                                                  .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                 (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata),   //                                                  .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest               (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                                  .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                                  .chipselect
		.led_pio_s1_address                                      (mm_interconnect_1_led_pio_s1_address),                        //                                        led_pio_s1.address
		.led_pio_s1_write                                        (mm_interconnect_1_led_pio_s1_write),                          //                                                  .write
		.led_pio_s1_readdata                                     (mm_interconnect_1_led_pio_s1_readdata),                       //                                                  .readdata
		.led_pio_s1_writedata                                    (mm_interconnect_1_led_pio_s1_writedata),                      //                                                  .writedata
		.led_pio_s1_chipselect                                   (mm_interconnect_1_led_pio_s1_chipselect),                     //                                                  .chipselect
		.sysid_control_slave_address                             (mm_interconnect_1_sysid_control_slave_address),               //                               sysid_control_slave.address
		.sysid_control_slave_readdata                            (mm_interconnect_1_sysid_control_slave_readdata),              //                                                  .readdata
		.timer_0_s1_address                                      (mm_interconnect_1_timer_0_s1_address),                        //                                        timer_0_s1.address
		.timer_0_s1_write                                        (mm_interconnect_1_timer_0_s1_write),                          //                                                  .write
		.timer_0_s1_readdata                                     (mm_interconnect_1_timer_0_s1_readdata),                       //                                                  .readdata
		.timer_0_s1_writedata                                    (mm_interconnect_1_timer_0_s1_writedata),                      //                                                  .writedata
		.timer_0_s1_chipselect                                   (mm_interconnect_1_timer_0_s1_chipselect)                      //                                                  .chipselect
	);

	nios2_control_irq_mapper irq_mapper (
		.clk           (altpll_0_c0_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_cpu_irq_irq)               //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_0_c1_clk),                    //       receiver_clk.clk
		.sender_clk     (altpll_0_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (altpll_0_c1_clk),                    //       receiver_clk.clk
		.sender_clk     (altpll_0_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (altpll_0_c1_clk),                    //       receiver_clk.clk
		.sender_clk     (altpll_0_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (nios2_cpu_debug_reset_request_reset), // reset_in1.reset
		.clk            (altpll_0_c0_clk),                     //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (nios2_cpu_debug_reset_request_reset), // reset_in1.reset
		.clk            (altpll_0_c1_clk),                     //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
